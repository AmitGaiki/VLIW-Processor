module mux2to1_23b(input enable, input [22:0] in1,input [22:0] in2, input sel,output reg[22:0] tagOut); 
   
 always @( in1,in2, sel,enable)
  
    if(enable) 
      begin
      case (sel)
      1'b0 : tagOut= in1;
      1'b1 : tagOut= in2;
      endcase
      end
    else tagOut = 23'd0;

endmodule

module mux2to1_64b(input enable, input [63:0] in1,input [63:0] in2, input sel,output reg[63:0] tagOut); 
   
 always @( in1,in2, sel,enable)
  
    if(enable) 
      begin
      case (sel)
      1'b0 : tagOut= in1;
      1'b1 : tagOut= in2;
      endcase
      end
    else tagOut = 64'd0;

endmodule

module mux2to1_22b(input enable, input [21:0] in1,input [21:0] in2, input sel,output reg[21:0] tagOut); 
   
 always @( in1,in2, sel,enable)
  
    if(enable) 
      begin
      case (sel)
      1'b0 : tagOut= in1;
      1'b1 : tagOut= in2;
      endcase
      end
    else tagOut = 22'd0;

endmodule

module mux8to1_8b(input enable, input [7:0] in0,in1,in2,in3,in4,in5,in6,in7,input [2:0] sel,output reg[7:0] out);
  always @(enable, in0,in1,in2,in3,in4,in5,in6,in7,sel)
  if(enable) begin
  case(sel)
    3'b000 : out = in0;
    3'b001 : out = in1;
    3'b010 : out = in2;
    3'b011 : out = in3;
    3'b100 : out = in4;
    3'b101 : out = in5;
    3'b110 : out = in6;
    3'b111 : out = in7;
  endcase
  end
endmodule

module mux64to1_23b(input enable, input[22:0] in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,
  in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,
  in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,
  in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,
  in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,
  in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,
  in60,in61,in62,in63,
    input [5:0] sel,output reg[22:0] out);
  always @(enable, in0,in1,in2,in3,in4,in5,in6,in7,in9,
          in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,
          in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,
          in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,
          in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,
          in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,
          in60,in61,in62,in63,sel)
  if(enable) begin
  case(sel)
    6'b000000 : out = in0;
    6'b000001 : out = in1;
    6'b000010 : out = in2;
    6'b000011 : out = in3;
    6'b000100 : out = in4;
    6'b000101 : out = in5;
    6'b000110 : out = in6;
    6'b000111 : out = in7;
	6'b001000 : out = in8;
    6'b001001 : out = in9;
    6'b001010 : out = in10;
    6'b001011 : out = in11;
    6'b001100 : out = in12;
    6'b001101 : out = in13;
    6'b001110 : out = in14;
    6'b001111 : out = in15;
	6'b010000 : out = in16;
    6'b010001 : out = in17;
    6'b010010 : out = in18;
    6'b010011 : out = in19;
    6'b010100 : out = in20;
    6'b010101 : out = in21;
    6'b010110 : out = in22;
    6'b010111 : out = in23;
	6'b011000 : out = in24;
    6'b011001 : out = in25;
    6'b011010 : out = in26;
    6'b011011 : out = in27;
    6'b011100 : out = in28;
    6'b011101 : out = in29;
    6'b011110 : out = in30;
    6'b011111 : out = in31;
	6'b100000 : out = in32;
    6'b100001 : out = in33;
    6'b100010 : out = in34;
    6'b100011 : out = in35;
    6'b100100 : out = in36;
    6'b100101 : out = in37;
    6'b100110 : out = in38;
    6'b100111 : out = in39;
	6'b101000 : out = in40;
    6'b101001 : out = in41;
    6'b101010 : out = in42;
    6'b101011 : out = in43;
    6'b101100 : out = in44;
    6'b101101 : out = in45;
    6'b101110 : out = in46;
    6'b101111 : out = in47;
	6'b110000 : out = in48;
    6'b110001 : out = in49;
    6'b110010 : out = in50;
    6'b110011 : out = in51;
    6'b110100 : out = in52;
    6'b110101 : out = in53;
    6'b110110 : out = in54;
    6'b110111 : out = in55;
	6'b111000 : out = in56;
    6'b111001 : out = in57;
    6'b111010 : out = in58;
    6'b111011 : out = in59;
    6'b111100 : out = in60;
    6'b111101 : out = in61;
    6'b111110 : out = in62;
    6'b111111 : out = in63;
  endcase
  end
  
endmodule

module mux64to1_64b(input enable, input[63:0] in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,
  in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,
  in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,
  in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,
  in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,
  in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,
  in60,in61,in62,in63,
    input [5:0] sel,output reg[63:0] out);
  always @(enable, in0,in1,in2,in3,in4,in5,in6,in7,in9,
          in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,
          in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,
          in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,
          in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,
          in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,
          in60,in61,in62,in63,sel)
  if(enable) begin
  case(sel)
    6'b000000 : out = in0;
    6'b000001 : out = in1;
    6'b000010 : out = in2;
    6'b000011 : out = in3;
    6'b000100 : out = in4;
    6'b000101 : out = in5;
    6'b000110 : out = in6;
    6'b000111 : out = in7;
	6'b001000 : out = in8;
    6'b001001 : out = in9;
    6'b001010 : out = in10;
    6'b001011 : out = in11;
    6'b001100 : out = in12;
    6'b001101 : out = in13;
    6'b001110 : out = in14;
    6'b001111 : out = in15;
	6'b010000 : out = in16;
    6'b010001 : out = in17;
    6'b010010 : out = in18;
    6'b010011 : out = in19;
    6'b010100 : out = in20;
    6'b010101 : out = in21;
    6'b010110 : out = in22;
    6'b010111 : out = in23;
	6'b011000 : out = in24;
    6'b011001 : out = in25;
    6'b011010 : out = in26;
    6'b011011 : out = in27;
    6'b011100 : out = in28;
    6'b011101 : out = in29;
    6'b011110 : out = in30;
    6'b011111 : out = in31;
	6'b100000 : out = in32;
    6'b100001 : out = in33;
    6'b100010 : out = in34;
    6'b100011 : out = in35;
    6'b100100 : out = in36;
    6'b100101 : out = in37;
    6'b100110 : out = in38;
    6'b100111 : out = in39;
	6'b101000 : out = in40;
    6'b101001 : out = in41;
    6'b101010 : out = in42;
    6'b101011 : out = in43;
    6'b101100 : out = in44;
    6'b101101 : out = in45;
    6'b101110 : out = in46;
    6'b101111 : out = in47;
	6'b110000 : out = in48;
    6'b110001 : out = in49;
    6'b110010 : out = in50;
    6'b110011 : out = in51;
    6'b110100 : out = in52;
    6'b110101 : out = in53;
    6'b110110 : out = in54;
    6'b110111 : out = in55;
	6'b111000 : out = in56;
    6'b111001 : out = in57;
    6'b111010 : out = in58;
    6'b111011 : out = in59;
    6'b111100 : out = in60;
    6'b111101 : out = in61;
    6'b111110 : out = in62;
    6'b111111 : out = in63;
  endcase
  end
  
endmodule

module mux64to1_1b(input enable, input in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,
    in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,
    in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,
    in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,
    in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,
    in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,
    in60,in61,in62,in63,
input [5:0] sel,output reg out);
  always @(enable, in0,in1,in2,in3,in4,in5,in6,in7,in9,
    in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,
    in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,
    in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,
    in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,
    in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,
    in60,in61,in62,in63,sel)
  if(enable) begin
  case(sel)
    6'b000000 : out = in0;
    6'b000001 : out = in1;
    6'b000010 : out = in2;
    6'b000011 : out = in3;
    6'b000100 : out = in4;
    6'b000101 : out = in5;
    6'b000110 : out = in6;
    6'b000111 : out = in7;
	6'b001000 : out = in8;
    6'b001001 : out = in9;
    6'b001010 : out = in10;
    6'b001011 : out = in11;
    6'b001100 : out = in12;
    6'b001101 : out = in13;
    6'b001110 : out = in14;
    6'b001111 : out = in15;
	6'b010000 : out = in16;
    6'b010001 : out = in17;
    6'b010010 : out = in18;
    6'b010011 : out = in19;
    6'b010100 : out = in20;
    6'b010101 : out = in21;
    6'b010110 : out = in22;
    6'b010111 : out = in23;
	6'b011000 : out = in24;
    6'b011001 : out = in25;
    6'b011010 : out = in26;
    6'b011011 : out = in27;
    6'b011100 : out = in28;
    6'b011101 : out = in29;
    6'b011110 : out = in30;
    6'b011111 : out = in31;
	6'b100000 : out = in32;
    6'b100001 : out = in33;
    6'b100010 : out = in34;
    6'b100011 : out = in35;
    6'b100100 : out = in36;
    6'b100101 : out = in37;
    6'b100110 : out = in38;
    6'b100111 : out = in39;
	6'b101000 : out = in40;
    6'b101001 : out = in41;
    6'b101010 : out = in42;
    6'b101011 : out = in43;
    6'b101100 : out = in44;
    6'b101101 : out = in45;
    6'b101110 : out = in46;
    6'b101111 : out = in47;
	6'b110000 : out = in48;
    6'b110001 : out = in49;
    6'b110010 : out = in50;
    6'b110011 : out = in51;
    6'b110100 : out = in52;
    6'b110101 : out = in53;
    6'b110110 : out = in54;
    6'b110111 : out = in55;
	6'b111000 : out = in56;
    6'b111001 : out = in57;
    6'b111010 : out = in58;
    6'b111011 : out = in59;
    6'b111100 : out = in60;
    6'b111101 : out = in61;
    6'b111110 : out = in62;
    6'b111111 : out = in63;	
  endcase
  end
endmodule

module decoder6to64(input [5:0] destReg, output reg [63:0] decOut);
always @(destReg)
  begin
    case(destReg)
      0: decOut =  64'b0000000000000000000000000000000000000000000000000000000000000001; 
      1: decOut =  64'b0000000000000000000000000000000000000000000000000000000000000010;
      2: decOut =  64'b0000000000000000000000000000000000000000000000000000000000000100;
      3: decOut =  64'b0000000000000000000000000000000000000000000000000000000000001000; 
      4: decOut =  64'b0000000000000000000000000000000000000000000000000000000000010000;
      5: decOut =  64'b0000000000000000000000000000000000000000000000000000000000100000;
      6: decOut =  64'b0000000000000000000000000000000000000000000000000000000001000000;
      7: decOut =  64'b0000000000000000000000000000000000000000000000000000000010000000;
      8: decOut =  64'b0000000000000000000000000000000000000000000000000000000100000000;
      9: decOut =  64'b0000000000000000000000000000000000000000000000000000001000000000;
      10: decOut = 64'b0000000000000000000000000000000000000000000000000000010000000000;
      11: decOut = 64'b0000000000000000000000000000000000000000000000000000100000000000;
      12: decOut = 64'b0000000000000000000000000000000000000000000000000001000000000000;
      13: decOut = 64'b0000000000000000000000000000000000000000000000000010000000000000;
      14: decOut = 64'b0000000000000000000000000000000000000000000000000100000000000000;
      15: decOut = 64'b0000000000000000000000000000000000000000000000001000000000000000;
      16: decOut = 64'b0000000000000000000000000000000000000000000000010000000000000000;
      17: decOut = 64'b0000000000000000000000000000000000000000000000100000000000000000;
      18: decOut = 64'b0000000000000000000000000000000000000000000001000000000000000000;
      19: decOut = 64'b0000000000000000000000000000000000000000000010000000000000000000;
      20: decOut = 64'b0000000000000000000000000000000000000000000100000000000000000000;
      21: decOut = 64'b0000000000000000000000000000000000000000001000000000000000000000;
      22: decOut = 64'b0000000000000000000000000000000000000000010000000000000000000000;
      23: decOut = 64'b0000000000000000000000000000000000000000100000000000000000000000;
      24: decOut = 64'b0000000000000000000000000000000000000001000000000000000000000000;
      25: decOut = 64'b0000000000000000000000000000000000000010000000000000000000000000;
      26: decOut = 64'b0000000000000000000000000000000000000100000000000000000000000000;
      27: decOut = 64'b0000000000000000000000000000000000001000000000000000000000000000;
      28: decOut = 64'b0000000000000000000000000000000000010000000000000000000000000000;
      29: decOut = 64'b0000000000000000000000000000000000100000000000000000000000000000;
      30: decOut = 64'b0000000000000000000000000000000001000000000000000000000000000000;
      31: decOut = 64'b0000000000000000000000000000000010000000000000000000000000000000;
      32: decOut = 64'b0000000000000000000000000000000100000000000000000000000000000000;
      33: decOut = 64'b0000000000000000000000000000001000000000000000000000000000000000;
      34: decOut = 64'b0000000000000000000000000000010000000000000000000000000000000000;
      35: decOut = 64'b0000000000000000000000000000100000000000000000000000000000000000;
      36: decOut = 64'b0000000000000000000000000001000000000000000000000000000000000000;
      37: decOut = 64'b0000000000000000000000000010000000000000000000000000000000000000;
      38: decOut = 64'b0000000000000000000000000100000000000000000000000000000000000000;
      39: decOut = 64'b0000000000000000000000001000000000000000000000000000000000000000;
      40: decOut = 64'b0000000000000000000000010000000000000000000000000000000000000000;
      41: decOut = 64'b0000000000000000000000100000000000000000000000000000000000000000;
      42: decOut = 64'b0000000000000000000001000000000000000000000000000000000000000000;
      43: decOut = 64'b0000000000000000000010000000000000000000000000000000000000000000;
      44: decOut = 64'b0000000000000000000100000000000000000000000000000000000000000000;
      45: decOut = 64'b0000000000000000001000000000000000000000000000000000000000000000;
      46: decOut = 64'b0000000000000000010000000000000000000000000000000000000000000000;
      47: decOut = 64'b0000000000000000100000000000000000000000000000000000000000000000;
      48: decOut = 64'b0000000000000001000000000000000000000000000000000000000000000000;
      49: decOut = 64'b0000000000000010000000000000000000000000000000000000000000000000;
      50: decOut = 64'b0000000000000100000000000000000000000000000000000000000000000000;
      51: decOut = 64'b0000000000001000000000000000000000000000000000000000000000000000;
      52: decOut = 64'b0000000000010000000000000000000000000000000000000000000000000000;
      53: decOut = 64'b0000000000100000000000000000000000000000000000000000000000000000;
      54: decOut = 64'b0000000001000000000000000000000000000000000000000000000000000000;
      55: decOut = 64'b0000000010000000000000000000000000000000000000000000000000000000;
      56: decOut = 64'b0000000100000000000000000000000000000000000000000000000000000000;
      57: decOut = 64'b0000001000000000000000000000000000000000000000000000000000000000;
      58: decOut = 64'b0000010000000000000000000000000000000000000000000000000000000000;
      59: decOut = 64'b0000100000000000000000000000000000000000000000000000000000000000;
      60: decOut = 64'b0001000000000000000000000000000000000000000000000000000000000000;
      61: decOut = 64'b0010000000000000000000000000000000000000000000000000000000000000;
      62: decOut = 64'b0100000000000000000000000000000000000000000000000000000000000000;
      63: decOut = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    endcase
  end                
endmodule

module comparator(input [22:0] in1, input [22:0] in2,output reg compOut);
  always@(in1, in2)
    begin
      if(in1 == in2)
        compOut = 1'b1;
      else
        compOut = 1'b0;
    end
endmodule

module orGate(input in1, input in2, output reg orOut);
  always@(in1, in2)
  begin
    if(in1 == 1 | in2 == 1)
      orOut = 1'b1;
    else
      orOut = 1'b0;
  end
endmodule